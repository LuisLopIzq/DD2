-- esto es un ejemplo que voy a comentar